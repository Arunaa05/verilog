module not_gate(input a,output c);
  assign c=~a;
endmodule
