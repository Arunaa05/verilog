module and_gate(input a,b,output c);
  assign c=a&b;
endmodule
